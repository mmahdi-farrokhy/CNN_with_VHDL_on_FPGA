library IEEE;
use IEEE.STD_LOGIC_1164.all;

package my_pkg is

end my_pkg;

package body my_pkg is

  type array8 is array (natural range <>) of std_logic_vector(7 downto 0);
 
end my_pkg;
